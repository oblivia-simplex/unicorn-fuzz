annel_stop_listening PKCS7_RECIP_INFO_it __GI_wcrtomb CMS_RecipientInfo_get0_pkey_ctx CRYPTO_dbg_get_options ECDH_get_default_method d2i_PBE2PARAM inflateInit2_ inflate_copyright mm_request_receive_expect d2i_PKCS7 platform_pre_fork CRYPTO_THREADID_set_callback OPENSSL_uni2asc __netlink_open _cs_write EC_POINT_is_on_curve UI_get_string_type X509_CRL_INFO_new BN_version RSA_set_default_method use_privsep BN_pseudo_rand X509_CRL_free EVP_PKEY_asn1_get0 zlibCompileFlags d2i_PKCS7_SIGN_ENVELOPE __GI_getuid PKCS7_set_signed_attributes a2i_ASN1_STRING s2i_ASN1_OCTET_STRING ECPARAMETERS_it RC4_options ERR_get_error_line_data BIO_ctrl_wpending BIO_f_asn1 ENGINE_get_default_RSA X509_get1_email DSA_up_ref ec_GFp_simple_field_sqr EVP_CIPHER_CTX_copy cms_SignerIdentifier_get0_signer_id EVP_PKEY_CTX_set_app_data SXNET_get_id_asc engine_table_doall BN_usub memset PKCS7_add_attrib_content_type i2d_PKCS7_bio sshkey_type_from_name ssh_packet_send EC_GROUP_get_curve_GFp fstatfs64 DES_decrypt3 MDC2_Final ENGINE_get_default_RAND DSO_load EC_KEY_get0_private_key setgid EVP_camellia_256_ecb __GI___sigaddset freeifaddrs __GI___ctype_b_loc i2d_PKCS8PrivateKey_nid_fp unlink BN_consttime_swap ERR_lib_error_string closefrom NCONF_default ec_pkey_meth putenv EVP_seed_ecb RSA_PSS_PARAMS_new EVP_CIPHER_CTX_flags ASN1_UNIVERSALSTRING_to_string _stdio_openlist_dec_use EVP_des_ede_ecb channel_after_select ISSUING_DIST_POINT_it strlcpy policy_data_new mm_key_sign RC2_ecb_encrypt BN_mod_sub ssh_packet_connection_af RSA_setup_blinding PEM_bytes_read_bio v3_idp d2i_PKCS12_fp __GI_mmap i2d_PROXY_CERT_INFO_EXTENSION PKCS12_MAC_DATA_free ENGINE_register_all_pkey_asn1_meths X509_CRL_sign active_state ECDSA_do_sign_ex __GI_strlcpy X509_policy_tree_level_count do_log2 syslogin_write_entry BN_mod_exp2_mont X509_ALGOR_dup BN_div EVP_CIPHER_CTX_set_padding d2i_X509_CERT_AUX a2d_ASN1_OBJECT asn1_set_choice_selector attrib_clear PKCS1_MGF1 __atexit_lock __GI_fread_unlocked CMS_signed_get_attr_by_OBJ crypto_sign_ed25519_ref_double_scalarmult_vartime _dl_pagesize OCSP_BASICRESP_new d2i_CRL_DIST_POINTS sshkey_ec_validate_private X509_signature_print PKCS7_add_signed_attribute EVP_PKEY_meth_set_derive CMS_get1_certs CRYPTO_ccm128_encrypt_ccm64 fakepw sshd_hostkey_sign X509_NAME_oneline ssh_hmac_init ASN1_TYPE_set_octetstring sshkey_equal_public sshkey_load_public UTF8_putc zlibVersion crypto_sign_ed25519_ref_sc25519_to32bytes POLICYQUALINFO_it fopencookie cms_RecipientInfo_kari_encrypt CRYPTO_THREADID_cpy mm_terminate PEM_write BIO_vprintf closelog CRYPTO_THREADID_set_numeric RSA_get_ex_new_index ec_GFp_simple_make_affine ASN1_item_d2i_fp asn1_GetSequence BN_generate_prime_ex v3_bcons ssh_krl_file_contains_key UI_add_verify_string i2d_ECPKParameters RAND_egd_bytes ASN1_STRING_free ECDSA_set_ex_data deflateReset PKCS12_key_gen_asc RSA_generate_key_ex DSA_sign_setup auth_request_forwarding PEM_write_PUBKEY check_defer lh_num_items Blowfish_decipher OBJ_NAME_cleanup ASN1_item_ex_free PKCS7_dataFinal X509_it X509_STORE_CTX_get_chain BF_options ec_GFp_simple_group_get_degree __GI_setresgid auth_rhosts_rsa_key_allowed BN_mod_sqr CONF_dump_fp cleanhostname EVP_aes_192_cfb8 ENGINE_set_default_ECDH d2i_RSAPublicKey_bio sigx_app ssh_digest_blocksize NCONF_new Camellia_EncryptBlock X509_STORE_CTX_purpose_inherit EC_KEY_set_group EVP_aes_192_cfb128 v3_ocsp_crlid __time_localtime_tzi X509_CRL_get0_by_cert d2i_ASN1_NULL __GI_strtoul i2d_ASN1_GENERALIZEDTIME ftello cms_EncryptedContent_init_bio d2i_PKCS12_MAC_DATA sshbuf_put_bignum1 BIO_f_cipher i2d_RSAPrivateKey_fp sshkey_ssh_name PKCS7_ENVELOPE_it ssh_packet_put_ecpoint EC_GROUP_get_seed_len PEM_write_RSAPrivateKey ENGINE_get_static_state EC_EX_DATA_clear_free_all_data sk_dup d2i_GENERAL_NAME ASN1_PCTX_new ENGINE_set_default_RSA i2d_ASN1_BOOLEAN __GI_fgets i2d_X509_VAL _CONF_new_data d2i_EXTENDED_KEY_USAGE X509_get_default_cert_file_env BN_get_word __pthread_mutex_unlock EVP_sha224 POLICY_MAPPING_new ASN1_ENUMERATED_new CMS_ContentInfo_free CRYPTO_memcmp i2a_ASN1_OBJECT OCSP_CERTSTATUS_new int_rsa_verify EC_POINT_make_affine crypto_si